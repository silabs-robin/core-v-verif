package uvm_pkg;
endpackage

`define  uvm_error(ID, MSG)  ;
`define  uvm_info(ID, MSG, VERBOSITY)  ;
`define  uvm_fatal(ID, MSG)  ;
